module buzzer_driver(
    input clk,
    input[4:0] note,
    output beep
    
)

endmodule